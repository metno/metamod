netcdf met_id_ch4 {
dimensions:
	data_status = 123 ;
variables:
	int data_status(data_status) ;
		data_status:units = "index" ;
		data_status:long_name = "Grid point status" ;
	float icedrift(data_status) ;
		icedrift:units = "km/24h" ;
		icedrift:long_name = "Ice displacement" ;
	float driftdirection(data_status) ;
		driftdirection:units = "degrees" ;
		driftdirection:long_name = "Displacement direction clock-wise from north" ;
	float correlation(data_status) ;
		correlation:units = "-" ;
		correlation:long_name = "Correlation coefficient" ;
	float latitude_reference(data_status) ;
		latitude_reference:units = "degrees_north" ;
		latitude_reference:long_name = "Latitude at start time" ;
	float longitude_reference(data_status) ;
		longitude_reference:units = "degrees_east" ;
		longitude_reference:long_name = "Longitude at start time" ;
	float latitude_compare(data_status) ;
		latitude_compare:units = "degrees_north" ;
		latitude_compare:long_name = "Latitude at stop time" ;
	float longitude_compare(data_status) ;
		longitude_compare:units = "degrees_east" ;
		longitude_compare:long_name = "Longitude at stop time" ;

// global attributes:
		:title = "METAMOD2 test data: Ice drift in Greenland seas" ;
		:abstract = "A 9 month ice drift data set based on VIS and IR data" ;
		:topiccategory = "Oceans" ;
		:keywords = "Ice drift, Arctic, IR, VIS, AVHRR, MCC" ;
		:activity_type = "Space borne instrument" ;
		:Conventions = "CF-1.0" ;
		:product_name = "Ice drift" ;
		:history = "2007-10-21 19:30:00 UTC creation" ;
		:area = "Arctic Ocean" ;
		:PI_name = "N.N" ;
		:contact = "n.n@nowhere.com ;
		:distribution_statement = "Free" ;
		:project_name = "METAMOD" ;
		:institution = "Some Meteorological Institute" ;
		:method = "Maximum Cross Correlation (MCC)" ;
		:correlation_window = "31x31 pixels" ;
		:original_data_desolution = "1000 m" ;
		:satelliteID_reference = "noaa17" ;
		:satelliteID_compare = "noaa17" ;
		:start_date = "2005-12-20 23:01:00 UTC" ;
		:stop_date = "2005-12-21 12:43:00 UTC" ;
		:platform = "AVHRR" ;
		:channel = 4 ;
		:northernsmost_latitude = 87.13695f ;
		:easternmost_longitude = 40.38439f ;
		:southernmost_latitude = 65.70739f ;
		:westernmost_longitude = -113.1208f ;
		:grid_spacing = 20 ;
		:leap_days = 0.5708333f ;
data:

 data_status = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0 ;

 icedrift = 18.86773, 12.63259, 25.08231, 16.15103, 10.65593, 18.62215, 
    19.97388, 24.77454, 24.77454, 7.222959, 6.316294, 8.759124, 22.77372, 
    10.51095, 11.7516, 11.7516, 10.21481, 17.86518, 12.63259, 7.432363, 
    24.52555, 18.62215, 23.56839, 18.03614, 23.56839, 13.3415, 15.6688, 
    11.7516, 13.3415, 11.7516, 11.7516, 10.21481, 10.21481, 12.63259, 
    11.21715, 12.63259, 21.0219, 10.21481, 12.63259, 12.63259, 10.21481, 
    22.4343, 11.7516, 12.63259, 12.63259, 10.21481, 12.63259, 10.21481, 
    18.62215, 12.63259, 12.63259, 10.21481, 11.7516, 10.21481, 8.759124, 
    24.33713, 22.4343, 9.909818, 14.12366, 11.21715, 14.12366, 8.759124, 
    9.909818, 12.63259, 12.63259, 12.63259, 8.759124, 9.909818, 9.909818, 
    8.759124, 21.16738, 15.06977, 9.909818, 9.909818, 8.759124, 11.21715, 
    8.759124, 10.21481, 12.38727, 11.21715, 10.21481, 10.21481, 11.21715, 
    11.07951, 8.759124, 11.21715, 11.21715, 11.21715, 12.38727, 23.82739, 
    11.21715, 9.909818, 10.21481, 11.21715, 12.63259, 8.759124, 10.21481, 
    11.21715, 8.759124, 10.21481, 9.909818, 9.909818, 14.86473, 14.86473, 
    16.52668, 14.44592, 17.25347, 23.04166, 8.932589, 25.08231, 12.63259, 
    19.27007, 19.586, 21.9503, 22.77372, 13.3415, 17.60562, 1.751825, 
    18.94888, 10.51095, 12.63259, 12.38727, 12.63259 ;

 driftdirection = 107, 51, 177, 190, 213, 250, 331, 308, 253, 197, 188, 190, 
    331, 241, 204, 201, 199, 157, 201, 192, 59, 282, 188, 213, 25, 203, 201, 
    213, 204, 204, 205, 202, 204, 203, 200, 207, 14, 200, 201, 203, 207, 205, 
    219, 199, 204, 204, 205, 229, 8, 203, 204, 208, 216, 225, 225, 115, 5, 
    191, 207, 200, 212, 228, 222, 202, 203, 204, 228, 222, 224, 218, 79, 201, 
    222, 224, 218, 222, 314, 348, 195, 216, 210, 212, 221, 210, 212, 229, 
    218, 224, 219, 117, 219, 214, 225, 219, 226, 220, 227, 221, 217, 225, 
    212, 214, 211, 213, 277, 323, 152, 318, 230, 296, 159, 307, 19, 324, 3, 
    228, 121, 197, 51, 191, 225, 198, 224 ;

 correlation = 0.7228356, 0.6985091, 0.6895878, 0.8370177, 0.7414688, 
    0.7261565, 0.7850716, 0.6726226, 0.7026024, 0.6729978, 0.7434388, 
    0.6228983, 0.628437, 0.6968202, 0.7501463, 0.6071896, 0.6073906, 
    0.7678297, 0.6064097, 0.7184624, 0.7491828, 0.662697, 0.6533465, 
    0.7227872, 0.690384, 0.7383977, 0.7439724, 0.6209559, 0.6018878, 
    0.6675799, 0.6484529, 0.6318137, 0.642721, 0.6532685, 0.6596028, 
    0.6786592, 0.6609755, 0.6251299, 0.7048455, 0.776201, 0.660484, 
    0.6055418, 0.683588, 0.7284984, 0.77238, 0.7573296, 0.7415259, 0.6416384, 
    0.732261, 0.6428371, 0.6960241, 0.7177382, 0.675419, 0.7279937, 
    0.6238618, 0.7196127, 0.641937, 0.6722608, 0.7757108, 0.6342916, 
    0.6637048, 0.6959035, 0.758478, 0.6904032, 0.7200257, 0.7235466, 
    0.7608003, 0.6947426, 0.6214306, 0.7109115, 0.7262788, 0.7229854, 
    0.6830812, 0.7231696, 0.7114668, 0.726337, 0.605737, 0.781488, 0.6383235, 
    0.6301147, 0.6471839, 0.7208334, 0.6567384, 0.8008388, 0.6548765, 
    0.6406285, 0.6254043, 0.6280909, 0.7264587, 0.6006162, 0.8386912, 
    0.6059786, 0.7344838, 0.797646, 0.6921596, 0.8065558, 0.73342, 0.7701963, 
    0.6191874, 0.7028933, 0.7139535, 0.6256088, 0.7329722, 0.8057995, 
    0.7282466, 0.8599357, 0.6515103, 0.6725773, 0.7779896, 0.660561, 
    0.8077152, 0.8333863, 0.6317897, 0.8784321, 0.7546195, 0.7401313, 
    0.6388226, 0.6453705, 0.7195215, 0.9444397, 0.871905, 0.9252692, 0.9281076 ;

 latitude_reference = 87.13695, 85.83435, 85.91528, 85.50426, 85.67426, 
    86.50255, 85.26269, 86.25087, 85.51595, 85.99805, 86.6302, 86.63315, 
    85.42647, 86.77427, 86.0967, 85.71577, 85.83692, 85.91391, 85.65726, 
    85.76065, 85.85841, 85.95013, 85.50522, 85.78747, 85.94452, 84.5479, 
    84.67429, 85.44725, 84.41398, 84.65703, 84.77306, 84.88509, 84.99284, 
    85.09604, 85.19438, 85.28757, 85.77245, 84.51424, 84.73607, 84.84069, 
    84.94077, 85.21091, 85.28996, 84.36904, 84.68652, 84.3287, 84.5305, 
    85.26648, 81.52092, 84.1765, 84.27676, 84.3728, 84.55124, 85.00891, 
    85.113, 81.56982, 81.26649, 83.92087, 84.02251, 84.12013, 84.30254, 
    84.95074, 84.96449, 83.6649, 83.76778, 83.86687, 84.76723, 84.7805, 
    84.78728, 84.78754, 83.40866, 83.51267, 84.59653, 84.60307, 84.60332, 
    84.59727, 82.47599, 82.08151, 83.55115, 84.41256, 84.41888, 84.41912, 
    84.41328, 84.29411, 84.21661, 84.2286, 84.23473, 83.8105, 83.8327, 
    81.43663, 83.53224, 83.5693, 83.31147, 83.35239, 83.38842, 83.1325, 
    83.17234, 83.20741, 82.86206, 82.90993, 82.95331, 82.99211, 82.55305, 
    82.59431, 79.30158, 78.27219, 78.24416, 78.01498, 77.98756, 77.84367, 
    78.02226, 77.80838, 75.04537, 72.37893, 71.25632, 71.24609, 71.17081, 
    67.60884, 67.43893, 65.88118, 65.84789, 65.73913, 65.70739 ;

 longitude_reference = 40.38439, 39.28407, -113.1208, -112.6912, -111.7634, 
    -105.788, -111.4736, -104.7027, -107.426, -103.7543, -92.8668, -88.42593, 
    -97.03241, -74.25042, -84.80431, -87.0169, -85.12958, -79.49555, 
    -80.12329, -78.08289, -75.94324, -73.70335, -78.76983, -72.49777, 
    -67.86726, -89.02847, -87.60123, -75.54683, -87.71323, -84.80465, 
    -83.25078, -81.62752, -79.93289, -78.16525, -76.32337, -74.40651, 
    -31.2102, -83.57103, -80.42933, -78.75954, -77.02209, -71.3981, 
    -69.38711, -82.4006, -77.65393, -79.78714, -76.61111, -55.19267, 
    11.71629, -78.75161, -77.2159, -75.62653, -72.28593, -58.98998, 
    -52.67992, 9.981476, 11.3691, -79.23119, -77.76921, -76.25758, -73.08423, 
    -50.32458, -48.23378, -79.67198, -78.27726, -76.8365, -50.13711, 
    -48.11953, -46.09419, -44.0661, -80.07845, -78.7453, -48.01308, 
    -46.05679, -44.09803, -42.14137, -0.7820017, 2.087021, -75.10748, 
    -47.91364, -46.02185, -44.12784, -42.23573, -32.94378, -49.64619, 
    -47.82055, -45.98916, -52.77478, -51.07669, -0.6868031, -57.41529, 
    -55.81023, -58.61858, -57.07354, -55.51048, -58.25631, -56.74984, 
    -55.22672, -60.79909, -59.3651, -57.91251, -56.44283, -58.66121, 
    -57.27497, -6.138511, -5.594735, -6.857034, -5.473473, -6.708872, 
    -7.246143, -9.87333, -8.459062, -16.02032, -20.12095, -19.26752, 
    -20.51789, -20.01103, -27.72596, -27.86345, -34.3638, -33.93948, 
    -34.86547, -34.443 ;

 latitude_compare = 87.10603, 85.87624, 85.78345, 85.4205, 85.62697, 
    86.46845, 85.35468, 86.33051, 85.4752, 85.96173, 86.59731, 86.58768, 
    85.53046, 86.74686, 86.03996, 85.65813, 85.78603, 85.82732, 85.59521, 
    85.72237, 85.92328, 85.97018, 85.38245, 85.70795, 86.05646, 84.48315, 
    84.59721, 85.39521, 84.34988, 84.60036, 84.71707, 84.83538, 84.94375, 
    85.03487, 85.1389, 85.22821, 85.8798, 84.46388, 84.67394, 84.77927, 
    84.89285, 85.10365, 85.24178, 84.30618, 84.62561, 84.2797, 84.47009, 
    85.23094, 81.61761, 84.11512, 84.21609, 84.32551, 84.50123, 84.97081, 
    85.08057, 81.51566, 81.3836, 83.8697, 83.95656, 84.06473, 84.23956, 
    84.91968, 84.92549, 83.60316, 83.70665, 83.80639, 84.7363, 84.74158, 
    84.7496, 84.75106, 83.42827, 83.43858, 84.55769, 84.56543, 84.56684, 
    84.55297, 82.50797, 82.13393, 83.48824, 84.36459, 84.37228, 84.37343, 
    84.36893, 84.24384, 84.1776, 84.18938, 84.18794, 83.76766, 83.78193, 
    81.37881, 83.48629, 83.52617, 83.2737, 83.30667, 83.342, 83.09714, 
    83.13583, 83.16292, 82.82545, 82.87169, 82.90917, 82.9487, 82.48631, 
    82.52856, 79.31155, 78.33264, 78.16454, 78.10438, 77.95732, 77.8997, 
    77.96082, 77.86791, 75.14153, 72.46968, 71.37311, 71.1999, 71.12451, 
    67.60035, 67.49956, 65.82903, 65.80257, 65.67978, 65.6617 ;

 longitude_compare = 42.26484, 39.99841, -113.0301, -112.872, -112.1606, 
    -107.2875, -112.0947, -106.2992, -109.0026, -103.914, -92.94906, 
    -88.55653, -97.78754, -75.10134, -85.1633, -87.31516, -85.36662, 
    -78.98683, -80.43607, -78.19116, -74.38586, -75.06515, -78.98997, 
    -73.19676, -67.10081, -89.31088, -87.91242, -75.965, -88.00397, 
    -85.06784, -83.53637, -81.855, -80.18182, -78.467, -76.56171, -74.76797, 
    -30.84317, -83.76566, -80.68439, -79.03952, -77.29619, -71.98112, 
    -69.85659, -82.61752, -77.93848, -80.00839, -76.89909, -55.67929, 
    11.80834, -79.00002, -77.48488, -75.8849, -72.66627, -59.42368, 
    -53.06279, 10.76676, 11.43789, -79.3223, -78.09457, -76.45335, -73.47806, 
    -50.70999, -48.62627, -79.89162, -78.51414, -77.09137, -50.51018, 
    -48.49912, -46.4891, -44.37472, -79.12366, -78.99034, -48.38058, 
    -46.43855, -44.39595, -42.5532, -1.034632, 2.005969, -75.25494, 
    -48.26445, -46.29517, -44.41674, -42.63334, -33.23841, -49.88818, 
    -48.25685, -46.34496, -53.14893, -51.45422, 0.0539666, -57.74162, 
    -56.06967, -58.94478, -57.39344, -55.9207, -58.50164, -57.07959, 
    -55.55206, -61.02233, -59.66889, -58.13638, -56.67709, -58.97144, 
    -57.59926, -6.600714, -5.816657, -6.651825, -5.861371, -6.878814, 
    -7.808252, -9.759259, -8.842967, -15.89358, -20.34419, -19.24764, 
    -20.67494, -19.771, -27.73288, -27.66878, -34.38768, -34.04886, 
    -34.91297, -34.55077 ;
}
